    ����          FAssembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null   SaveGameObj   BuyGj�System.Collections.Generic.List`1[[UnityEngine.GameObject, UnityEngine.CoreModule, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   	      MUnityEngine.CoreModule, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null   �System.Collections.Generic.List`1[[UnityEngine.GameObject, UnityEngine.CoreModule, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  UnityEngine.GameObject[]   	         